typedef enum logic [2:0] {
    FETCH = 3'b000,
    FETCH_IMEM = 3'b001,
    DECODE = 3'b010,
    EXECUTE = 3'b011,
    MEMORY = 3'b100,
    WRITEBACK = 3'b101,
    HALT = 3'b110
} cpu_state_t;

module Core(
    input clk,
    input rst,
    input [31:0] data_in,
    output logic [31:0] data_out,
    output logic [31:0] address,
    output logic write_enable,
    output logic [7:0] debug_out
);

    cpu_state_t state;

    (* ram_style = "distributed" *) logic [31:0] gp_registers[0:7];
    (* ram_style = "distributed" *) logic [31:0] special_registers[0:7];

    logic [3:0] rsrc1;
    logic [3:0] rsrc2;
    logic [3:0] rdest;

    logic [31:0] immediate;
    logic [31:0] imem;

    logic [7:0] opcode;
    control_signal_t control_signal;
    logic [3:0] alu_opcode;

    logic[31:0] rsrc1_value;
    logic[31:0] rsrc2_value;
    logic [31:0] alu_result;

    CU cu (
        .clk(clk),
        .rst(rst),
        .opcode(opcode),
        .control_signal(control_signal),
        .alu_opcode(alu_opcode)
    );

    ALU alu (
        .clk(clk),
        .opcode(alu_opcode),
        .a(rsrc1_value),
        .b(control_signal.alu_b_use_immediate ? immediate : rsrc2_value),
        .result(alu_result)
    );

    logic enable_jump;
    always_comb begin
        unique case (control_signal.jump_condition)
            JC_ALWAYS: enable_jump = 1'b1;
            JC_IF_ZERO: enable_jump = (rsrc1_value == 32'b0);
            JC_IF_NOT_ZERO: enable_jump = (rsrc1_value != 32'b0);
            JC_IF_NEGATIVE: enable_jump = rsrc1_value[31];
            JC_IF_NOT_NEGATIVE: enable_jump = ~rsrc1_value[31];
            default: enable_jump <= 1'b0; // Invalid state
        endcase
    end

    logic [31:0] ip_inc;
    always_comb begin
        unique case (data_in[7:5])
            3'b000: ip_inc = 1;
            3'b001: ip_inc = 2;
            3'b010: ip_inc = 1;
            3'b011: ip_inc = 2;
            3'b100: ip_inc = 2;
            3'b101: ip_inc = 3;
            3'b110: ip_inc = 2;
            default: ip_inc = 0; // Invalid state
        endcase
    end

    logic [31:0] ip_next;

    always_ff @(posedge clk or posedge rst) begin
        if (rst) begin
            state <= FETCH;
            address <= 32'b0;
            data_out <= 32'b0;
            debug_out <= 8'b11111111;

            for (integer i = 0; i < 8; i = i + 1) begin
                gp_registers[i] <= 32'b0;
                special_registers[i] <= 32'b0;
            end
        end else begin
            case (state)
                FETCH: begin
                    (* use_dsp = "yes" *) ip_next = special_registers[0] + ip_inc;
                    opcode <= data_in[7:0];
                    debug_out <= data_in[7:0];
                    case (data_in[7:5])
                        3'b000: begin // No extra values
                            state <= DECODE;
                        end
                        3'b001: begin // Immediate
                            // For now, assume 8 bits. This may change in the future
                            immediate <= {24'b0, data_in[15:8]};
                            state <= DECODE;
                        end
                        3'b010: begin // Address
                            address <= ip_next;
                            state <= FETCH_IMEM;
                        end
                        3'b011: begin // Immediate + Address
                            immediate <= {24'b0, data_in[15:8]};
                            address <= ip_next;
                            state <= FETCH_IMEM;
                        end
                        3'b100: begin // Register
                            rsrc1 <= data_in[15:12];
                            rsrc2 <= data_in[11:8];
                            // Let's assume that the first source is also the destination
                            rdest <= data_in[15:12];
                            state <= DECODE;
                        end
                        3'b101: begin // Register + Immediate
                            rsrc1 <= data_in[15:12];
                            rsrc2 <= data_in[11:8];
                            rdest <= data_in[15:12];
                            immediate <= {24'b0, data_in[23:16]};
                            state <= DECODE;
                        end
                        3'b110: begin // Register + Address
                            rsrc1 <= data_in[15:12];
                            rsrc2 <= data_in[11:8];
                            rdest <= data_in[15:12];
                            address <= ip_next;
                            state <= FETCH_IMEM;
                        end
                        3'b111: begin // Invalid state
                            state <= HALT;
                        end
                    endcase
                    special_registers[0] <= ip_next;
                end
                FETCH_IMEM: begin
                    debug_out <= 8'b00000010;
                    imem <= data_in;
                    special_registers[0] <= special_registers[0] + 4;
                    state <= DECODE;
                end
                DECODE: begin
                    debug_out <= 8'b00000011;
                    rsrc1_value = lookup_gp_register(rsrc1);
                    rsrc2_value = lookup_gp_register(rsrc2);
                    state <= EXECUTE;
                end
                EXECUTE: begin
                    debug_out <= 8'b00000100;
                    if (control_signal.halt) begin
                        state <= HALT;
                    end else begin
                        address <= imem;
                        state <= MEMORY;

                        if (enable_jump) begin
                            case (control_signal.jmp_src)
                                JS_NO_JUMP_SRC: begin end // No Jump
                                JS_JUMP_SRC_RDEST: special_registers[0] <= lookup_gp_register(rdest);
                                JS_JUMP_SRC_IMMEDIATE: special_registers[0] <= add_immediate_8(special_registers[0], immediate);
                                JS_JUMP_SRC_ADDR: special_registers[0] <= imem;
                                default: state <= HALT; // Invalid state
                            endcase
                        end
                    end
                end
                MEMORY: begin
                    debug_out <= 8'b00000101;
                    case (control_signal.write_memory_src)
                        WM_WRITE_SRC_RSRC1: begin
                            data_out <= lookup_gp_register(rsrc1);
                            write_enable <= 1'b1;
                        end
                        WM_WRITE_SRC_IMMEDIATE: begin
                            data_out <= immediate;
                            write_enable <= 1'b1;
                        end
                    endcase
                    state <= WRITEBACK;
                end
                WRITEBACK: begin;
                    debug_out <= 8'b00000110;
                    write_enable <= 1'b0;

                    case (control_signal.write_register_src)
                        WR_WRITE_SRC_RDEST: write_gp_register(rdest, alu_result);
                        WR_WRITE_SRC_RSRC2: write_gp_register(rdest, rsrc2_value);
                        WR_WRITE_SRC_MEMORY: write_gp_register(rdest, data_in);
                        WR_WRITE_SRC_IMMEDIATE: write_gp_register(rdest, immediate);
                    endcase

                    state <= FETCH;
                    address <= special_registers[0];
                end
                HALT: begin
                    debug_out <= 8'b11111111;
                end
            endcase
        end
    end

    task automatic write_gp_register;
        input [2:0] index;
        input [31:0] value;
        begin
            gp_registers[index] <= value;
        end
    endtask

    function [31:0] lookup_gp_register;
        input [2:0] index;
        begin
            lookup_gp_register = gp_registers[index];
        end
    endfunction

    function [31:0] add_immediate_8;
        input [31:0] value;
        input [31:0] immediate;
        logic [7:0] imm8;
        logic signed [31:0] sign_extended_imm;
        begin
            imm8 = immediate[7:0];
            sign_extended_imm = {{24{imm8[7]}}, imm8};
            (* use_dsp = "yes" *) add_immediate_8 = value + sign_extended_imm;
        end
    endfunction


endmodule